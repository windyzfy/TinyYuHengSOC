module regs(
          input wire clk,
          input wire rst_n,
          //from id
          input wire [4:0] reg1_raddr_i,
          input wire [4:0] reg2_raddr_i,
          //to id
          output reg [31:0] reg1_rdata_o,
          output reg [31:0] reg2_rdata_o
);
          reg [31:0] regs[0:31];        //定义寄存器组
          always @(*)begin
                    if(!rst_n)begin
                              reg1_rdata_o = 32'b0;
                    end
                    else if(reg1_raddr_i == 0)begin         //访问0号寄存器，值永远为0
                              reg1_rdata_o = 32'b0;
                    end
                    else begin
                              reg1_rdata_o = regs[reg1_raddr_i];
                    end
          end
          
          always @(*)begin
                    if(!rst_n)begin
                              reg2_rdata_o = 32'b0;
                    end
                    else if(reg2_raddr_i == 0)begin         //访问0号寄存器，值永远为0
                              reg2_rdata_o = 32'b0;
                    end
                    else begin
                              reg2_rdata_o = regs[reg2_raddr_i];
                    end
          end

endmodule